fb[30][14] <= 1'b0;
fb[30][16] <= 1'b0;
fb[29][12] <= 1'b0;
fb[29][18] <= 1'b0;
fb[28][10] <= 1'b0;
fb[28][20] <= 1'b0;
fb[26][9] <= 1'b0;
fb[26][21] <= 1'b0;
fb[24][8] <= 1'b0;
fb[24][22] <= 1'b0;
fb[22][8] <= 1'b0;
fb[22][22] <= 1'b0;
fb[20][9] <= 1'b0;
fb[20][21] <= 1'b0;
fb[18][10] <= 1'b0;
fb[18][20] <= 1'b0;
fb[17][12] <= 1'b0;
fb[17][18] <= 1'b0;
fb[16][14] <= 1'b0;
fb[16][16] <= 1'b0;
fb[6][10] <= 1'b0;
fb[6][11] <= 1'b0;
fb[6][12] <= 1'b0;
fb[6][13] <= 1'b0;
fb[6][14] <= 1'b0;
fb[6][16] <= 1'b0;
fb[6][17] <= 1'b0;
fb[6][18] <= 1'b0;
fb[6][19] <= 1'b0;
fb[6][20] <= 1'b0;
fb[5][10] <= 1'b0;
fb[5][14] <= 1'b0;
fb[5][20] <= 1'b0;
fb[4][10] <= 1'b0;
fb[4][14] <= 1'b0;
fb[4][20] <= 1'b0;
fb[3][10] <= 1'b0;
fb[3][14] <= 1'b0;
fb[3][20] <= 1'b0;
fb[2][10] <= 1'b0;
fb[2][14] <= 1'b0;
fb[2][20] <= 1'b0;
fb[1][10] <= 1'b0;
fb[1][14] <= 1'b0;
fb[1][20] <= 1'b0;
fb[0][10] <= 1'b0;
fb[0][11] <= 1'b0;
fb[0][12] <= 1'b0;
fb[0][13] <= 1'b0;
fb[0][14] <= 1'b0;
fb[0][20] <= 1'b0;
