fb[38][13] <= 1'b1;
fb[38][15] <= 1'b1;
fb[38][17] <= 1'b1;
fb[37][10] <= 1'b1;
fb[37][20] <= 1'b1;
fb[36][8] <= 1'b1;
fb[36][22] <= 1'b1;
fb[34][5] <= 1'b1;
fb[34][25] <= 1'b1;
fb[32][3] <= 1'b1;
fb[32][27] <= 1'b1;
fb[30][2] <= 1'b1;
fb[30][28] <= 1'b1;
fb[28][1] <= 1'b1;
fb[28][29] <= 1'b1;
fb[25][0] <= 1'b1;
fb[25][30] <= 1'b1;
fb[23][0] <= 1'b1;
fb[23][30] <= 1'b1;
fb[21][0] <= 1'b1;
fb[21][30] <= 1'b1;
fb[18][1] <= 1'b1;
fb[18][29] <= 1'b1;
fb[16][2] <= 1'b1;
fb[16][28] <= 1'b1;
fb[14][3] <= 1'b1;
fb[14][27] <= 1'b1;
fb[12][5] <= 1'b1;
fb[12][25] <= 1'b1;
fb[10][8] <= 1'b1;
fb[10][22] <= 1'b1;
fb[9][10] <= 1'b1;
fb[9][20] <= 1'b1;
fb[8][13] <= 1'b1;
fb[8][15] <= 1'b1;
fb[8][17] <= 1'b1;
fb[6][14] <= 1'b1;
fb[6][16] <= 1'b1;
fb[6][17] <= 1'b1;
fb[6][18] <= 1'b1;
fb[6][19] <= 1'b1;
fb[6][20] <= 1'b1;
fb[5][14] <= 1'b1;
fb[5][16] <= 1'b1;
fb[4][14] <= 1'b1;
fb[4][16] <= 1'b1;
fb[3][14] <= 1'b1;
fb[3][16] <= 1'b1;
fb[3][17] <= 1'b1;
fb[3][18] <= 1'b1;
fb[3][19] <= 1'b1;
fb[3][20] <= 1'b1;
fb[2][14] <= 1'b1;
fb[2][20] <= 1'b1;
fb[1][14] <= 1'b1;
fb[1][20] <= 1'b1;
fb[0][14] <= 1'b1;
fb[0][16] <= 1'b1;
fb[0][17] <= 1'b1;
fb[0][18] <= 1'b1;
fb[0][19] <= 1'b1;
fb[0][20] <= 1'b1;
