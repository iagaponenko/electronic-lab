fb[24][15] <= 1'b1;
fb[23][14] <= 1'b1;
fb[23][16] <= 1'b1;
fb[22][15] <= 1'b1;
fb[6][10] <= 1'b1;
fb[6][11] <= 1'b1;
fb[6][12] <= 1'b1;
fb[6][13] <= 1'b1;
fb[6][14] <= 1'b1;
fb[6][20] <= 1'b1;
fb[5][10] <= 1'b1;
fb[5][14] <= 1'b1;
fb[5][20] <= 1'b1;
fb[4][10] <= 1'b1;
fb[4][14] <= 1'b1;
fb[4][20] <= 1'b1;
fb[3][10] <= 1'b1;
fb[3][14] <= 1'b1;
fb[3][20] <= 1'b1;
fb[2][10] <= 1'b1;
fb[2][14] <= 1'b1;
fb[2][20] <= 1'b1;
fb[1][10] <= 1'b1;
fb[1][14] <= 1'b1;
fb[1][20] <= 1'b1;
fb[0][10] <= 1'b1;
fb[0][11] <= 1'b1;
fb[0][12] <= 1'b1;
fb[0][13] <= 1'b1;
fb[0][14] <= 1'b1;
fb[0][20] <= 1'b1;
