-- The rotary encoder which also includes a debouncer.

Library ieee;
Use ieee.std_logic_1164.All;
Use ieee.numeric_std.All;

Package rotary_encoder Is
End Package rotary_encoder;

Package Body rotary_encoder Is
End Package Body rotary_encoder;

