-- The frame buffer

Library ieee;
Use ieee.std_logic_1164.All;
Use ieee.numeric_std.All;

Package framebuffer Is
End Package framebuffer;

Package Body framebuffer Is
End Package Body framebuffer;

