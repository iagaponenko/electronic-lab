fb[33][14] <= 1'b0;
fb[33][16] <= 1'b0;
fb[32][11] <= 1'b0;
fb[32][19] <= 1'b0;
fb[31][9] <= 1'b0;
fb[31][21] <= 1'b0;
fb[30][8] <= 1'b0;
fb[30][22] <= 1'b0;
fb[29][7] <= 1'b0;
fb[29][23] <= 1'b0;
fb[27][6] <= 1'b0;
fb[27][24] <= 1'b0;
fb[24][5] <= 1'b0;
fb[24][25] <= 1'b0;
fb[22][5] <= 1'b0;
fb[22][25] <= 1'b0;
fb[19][6] <= 1'b0;
fb[19][24] <= 1'b0;
fb[17][7] <= 1'b0;
fb[17][23] <= 1'b0;
fb[16][8] <= 1'b0;
fb[16][22] <= 1'b0;
fb[15][9] <= 1'b0;
fb[15][21] <= 1'b0;
fb[14][11] <= 1'b0;
fb[14][19] <= 1'b0;
fb[13][14] <= 1'b0;
fb[13][16] <= 1'b0;
fb[6][14] <= 1'b0;
fb[6][16] <= 1'b0;
fb[6][17] <= 1'b0;
fb[6][18] <= 1'b0;
fb[6][19] <= 1'b0;
fb[6][20] <= 1'b0;
fb[5][14] <= 1'b0;
fb[5][16] <= 1'b0;
fb[5][20] <= 1'b0;
fb[4][14] <= 1'b0;
fb[4][16] <= 1'b0;
fb[4][20] <= 1'b0;
fb[3][14] <= 1'b0;
fb[3][16] <= 1'b0;
fb[3][20] <= 1'b0;
fb[2][14] <= 1'b0;
fb[2][16] <= 1'b0;
fb[2][20] <= 1'b0;
fb[1][14] <= 1'b0;
fb[1][16] <= 1'b0;
fb[1][20] <= 1'b0;
fb[0][14] <= 1'b0;
fb[0][16] <= 1'b0;
fb[0][17] <= 1'b0;
fb[0][18] <= 1'b0;
fb[0][19] <= 1'b0;
fb[0][20] <= 1'b0;
