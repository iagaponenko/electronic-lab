-- The dummy package. The package is required by the IDE for implementing
-- the SPI serializer(s).

Library ieee;
Use ieee.std_logic_1164.All;
Use ieee.numeric_std.All;

Package max7219 Is
End Package max7219;

Package Body max7219 Is
End Package Body max7219;

