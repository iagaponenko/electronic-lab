-- Implement an SPI-like serializer for MAX7219.
--
-- https://www.sparkfun.com/datasheets/Components/General/COM-09622-MAX7219-MAX7221.pdf

Library ieee;
Use ieee.std_logic_1164.All;
Use ieee.numeric_std.All;
Use ieee.math_real.All;

Entity spi_max7219 Is
    Port (
        -- Management interface
        rst      : In  std_logic;
        clk      : In  std_logic;
        start    : In  std_logic;
        data     : In  std_logic_vector(15 Downto 0);
        busy     : Out std_logic;
        -- SPI signals generated by the entity
        spi_clk  : Out std_logic;
        spi_load : Out std_logic;
        spi_din  : Out std_logic
    );
End Entity spi_max7219;


Architecture Behavioral Of spi_max7219 Is
    Type ProcessingState Is (IDLE, RUNNING);
    Signal state : ProcessingState := IDLE;
Begin
    bcd_compute_process : Process (clk, rst, start, state) Is
        Variable n : natural Range 0 To 15;
    Begin
        If rst Then
          	spi_clk  <= '0';
          	spi_load <= '0';
          	spi_din  <= 'X';
            state <= IDLE;
        ElsIf rising_edge(clk) Then
            Case state Is
                When IDLE =>
                    spi_load <= '0';
                    If start Then
                        state <= RUNNING;
                        n := 15;
                    	spi_clk  <= '1';
                        spi_din <= data(n);
                    End If;
                When RUNNING =>
                    spi_clk  <= '1';
                    If n = 0 Then
                    	spi_load <= '1';
                        state <= IDLE;
                    Else
                        n := n - 1;
                        spi_din <= data(n);
                    End If;
                When Others =>
                 	spi_clk  <= '0';
          	        spi_load <= '0';
                    spi_din <= 'X';
                    state <= IDLE;
            End Case;
        ElsIf falling_edge(clk) Then
            spi_clk  <= '0';
        End If;
    End Process bcd_compute_process;

    -- Device "busy" is set during when the last request is still being processed.
    -- The "start" command will be ignored in this state.
    busy <= '0' When state = IDLE    Else
            '1' When state = RUNNING Else
            'X';

End Architecture Behavioral;

