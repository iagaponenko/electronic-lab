fb[37][13] <= 1'b0;
fb[37][15] <= 1'b0;
fb[37][17] <= 1'b0;
fb[36][10] <= 1'b0;
fb[36][20] <= 1'b0;
fb[35][8] <= 1'b0;
fb[35][22] <= 1'b0;
fb[33][5] <= 1'b0;
fb[33][25] <= 1'b0;
fb[32][4] <= 1'b0;
fb[32][26] <= 1'b0;
fb[30][3] <= 1'b0;
fb[30][27] <= 1'b0;
fb[28][2] <= 1'b0;
fb[28][28] <= 1'b0;
fb[25][1] <= 1'b0;
fb[25][29] <= 1'b0;
fb[23][1] <= 1'b0;
fb[23][29] <= 1'b0;
fb[21][1] <= 1'b0;
fb[21][29] <= 1'b0;
fb[18][2] <= 1'b0;
fb[18][28] <= 1'b0;
fb[16][3] <= 1'b0;
fb[16][27] <= 1'b0;
fb[14][4] <= 1'b0;
fb[14][26] <= 1'b0;
fb[13][5] <= 1'b0;
fb[13][25] <= 1'b0;
fb[11][8] <= 1'b0;
fb[11][22] <= 1'b0;
fb[10][10] <= 1'b0;
fb[10][20] <= 1'b0;
fb[9][13] <= 1'b0;
fb[9][15] <= 1'b0;
fb[9][17] <= 1'b0;
fb[6][14] <= 1'b0;
fb[6][16] <= 1'b0;
fb[6][20] <= 1'b0;
fb[5][14] <= 1'b0;
fb[5][16] <= 1'b0;
fb[5][20] <= 1'b0;
fb[4][14] <= 1'b0;
fb[4][16] <= 1'b0;
fb[4][20] <= 1'b0;
fb[3][14] <= 1'b0;
fb[3][16] <= 1'b0;
fb[3][17] <= 1'b0;
fb[3][18] <= 1'b0;
fb[3][19] <= 1'b0;
fb[3][20] <= 1'b0;
fb[2][14] <= 1'b0;
fb[2][20] <= 1'b0;
fb[1][14] <= 1'b0;
fb[1][20] <= 1'b0;
fb[0][14] <= 1'b0;
fb[0][20] <= 1'b0;
