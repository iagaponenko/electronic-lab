-- A driver for the SPI-like serializer for MAX7219. The driver is meant
-- to be run on the Digilent Basys 3 development board.
--
-- 5 strips of 4 digits each, 20 digits in total
-- first strip is read, 4 strips are green
--
-- 4 rotary encoderers, of which 4 loqwer ones are used for incremending/decrementing
-- a value of the 4-decimal digit number by 1.

Library ieee;
Use ieee.std_logic_1164.All;
Use ieee.std_logic_unsigned.All;
Use ieee.numeric_std.All;
Use ieee.math_real.All;

Entity drive_spi_max7219_synt_20 Is
    Generic (
        NUM_RENCODERS : natural :=  5;
        NUM_SWITCHES  : natural := 16
    );
    Port (
        -- Input signals sent by the board into the module
        clk          : In  std_logic;   -- 100 MHz clock

        -- 5 push buttons on the FPGA board
        g_btn_up     : In  std_logic;
        g_btn_right  : In  std_logic;
        g_btn_down   : In  std_logic;
        g_btn_left   : In  std_logic;
        g_btn_center : In  std_logic;

        -- 16 control switches on the FPGA board
        g_sw         : In std_logic_vector(NUM_SWITCHES - 1 Downto 0);

        -- SPI signals generated by the entity. These are sent the output
        -- ports of the FPGA board.
        g_spi_clk    : Out std_logic;
        g_spi_load   : Out std_logic;
        g_spi_din    : Out std_logic;

        -- The clock that drives the serializer. It's sent to the output port
        -- of the FPGA board to allow external inspection and diagnostics.
        g_div_clk    : Out std_logic;

        -- Rotary encoder interface: channels 'a' and 'b', push button 'p'
        g_rencoder_a : In std_logic_vector(0 To NUM_RENCODERS - 1); 
        g_rencoder_b : In std_logic_vector(0 To NUM_RENCODERS - 1);
        g_rencoder_p : In std_logic_vector(0 To NUM_RENCODERS - 1);     -- pulled up

        -- Debug signals for the rotary encoder interface
        g_rencoder_left  : Out std_logic;
        g_rencoder_right : Out std_logic
     );
End Entity drive_spi_max7219_synt_20;

Architecture Rtl Of drive_spi_max7219_synt_20 Is

    -- Aliases for the inputs
    Alias rst_btn : std_logic Is g_btn_center;

    -- Using 4 out of 5.
    Constant DIGITS : natural := NUM_RENCODERS - 1;

    -- Key frequencies (Hz)
    Constant FREQ_CLK                  : natural := 100_000_000; 
    Constant FREQ_SPI_DRIVE_CLK        : natural :=   1_000_000;
    Constant FREQ_DISPLEY_UPDATE       : natural :=         500;
    Constant FREQ_RENCODER_CLK_PERIODS : natural :=     100_000;  -- corresponds to 10 ms minimum stable duration of the pressed button
    Constant FREQ_COUNTER_CLK          : natural :=          10;  -- counter for incrementing the number on the display

    Signal rst           : std_logic;
    Signal start         : std_logic;
    Signal busy          : std_logic;
    Signal spi_drive_clk : std_logic;
    Signal spi_load      : std_logic;
    Signal diag_state    : std_logic_vector(3 Downto 0);

    Constant HDR : std_logic_vector(3 Downto 0) := "0000";

    Subtype RegType  Is std_logic_vector(3 Downto 0);
    Subtype DataType Is std_logic_vector(7 Downto 0);

    Constant REG_NOP : RegType  := "0000";
    Constant D_NOP : DataType := "00000000";

    Constant NUM_STRIPS : natural := 5;
    Constant NUM_DIGITS_PER_STRIP : natural := 4;
    Constant NUM_DIGITS : natural := NUM_STRIPS * NUM_DIGITS_PER_STRIP;
    Subtype DataStreamType Is std_logic_vector(16 * NUM_DIGITS - 1  Downto 0);

    Constant NOP : DataStreamType :=
        HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP &
        HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP &
        HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP &
        HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP &
        HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP & HDR & REG_NOP & D_NOP;

    ---------------------
    -- Symbol matrixes --
    ---------------------

    Subtype SymbolMatrix Is std_logic_vector(63 Downto 0);
    Type DecimalNumbers Is Array (0 To 9) Of SymbolMatrix;
-- Very tiny: 3x5
--    Constant DECIMAL : DecimalNumbers := (
--          X"e0a0a0a0e0000000",
--          X"8080808080000000",
--          X"e020e080e0000000",
--          X"e080e080e0000000",
--          X"8080e0a0a0000000",
--          X"e080e020e0000000",
--          X"e0a0e020e0000000",
--          X"80808080e0000000",
--          X"e0a0e0a0e0000000",
--          X"e080e0a0e0000000"
--    );
--  Toll: 3x7
--    Constant DECIMAL : DecimalNumbers := (
--            X"e0a0a0a0a0a0e000",
--            X"8080808080808000",
--            X"e02020e08080e000",
--            X"e08080e08080e000",
--            X"808080e0a0a0a000",
--            X"e08080e02020e000",
--            X"e0a0a0e02020e000",
--            X"808080808080e000",
--            X"e0a0a0e0a0a0e000",
--            X"e08080e0a0a0e000"
--    );
--  Medimum: 4x7
    Constant DECIMAL : DecimalNumbers := (
            X"f09090909090f000",
            X"8080808080808000",
            X"f80808788080f800",
            X"f08080f08080f000",
            X"808080f090909000",
            X"f08080f01010f000",
            X"f09090f01010f000",
            X"808080808080f000",
            X"f09090f09090f000",
            X"f08080f09090f000"
    );
--  Medimum: 5x7
--    Constant DECIMAL : DecimalNumbers := (
--            X"f88888888888f800",
--            X"8080808080808000",
--            X"f80808f88080f800",
--            X"f88080f88080f800",
--            X"808080f888888800",
--            X"f88080f80808f800",
--            X"f88888f80808f800",
--            X"808080808080f800",
--            X"f88888f88888f800",
--            X"f88080f88888f800"
--    );
-- Very large: 7x8
--    Constant DECIMAL : DecimalNumbers := (
--        X"1c2222222222221c",
--        X"1c08080808080c08",
--        X"3e0408102020221c",
--        X"1c2220201820221c",
--        X"20203e2224283020",
--        X"1c2220201e02023e",
--        X"1c2222221e02221c",
--        X"040404081020203e",
--        X"1c2222221c22221c",
--        X"1c22203c2222221c"
--    );
    Subtype RowSelectorType Is natural Range 0 To 7;
    Function symbol_row(symbol : SymbolMatrix;
                        row_selector : RowSelectorType) Return DataType Is
        Constant IDX : natural Range 63 Downto 0 := (7 - row_selector) * 8;
    Begin
        Return symbol(IDX + 7 Downto IDX);
    End Function;

    Type RegRows Is Array (0 To 7) Of RegType;
    Constant REG_ROW  : RegRows := (
        "0001", "0010", "0011", "0100", "0101", "0110", "0111", "1000"
    );

    ---------------------------------------------------
    -- Set same data at the specified row of all digits
    ---------------------------------------------------
    Function set_row(row_selector : RowSelectorType;
                     data         : DataType) Return DataStreamType Is
        Variable result : DataStreamType;
        Variable pos_hdr_begin : integer;
        Variable pos_reg_begin : integer;
        Variable pos_dat_begin : integer;
    Begin
        For digit In NUM_DIGITS - 1 Downto 0 Loop
            pos_hdr_begin := (digit + 1) * 16 - 1;
            pos_reg_begin := pos_hdr_begin - 4;
            pos_dat_begin := pos_reg_begin - 4;
            result(pos_hdr_begin Downto pos_hdr_begin - 3) := HDR;
            result(pos_reg_begin Downto pos_reg_begin - 3) := REG_ROW(row_selector);
            result(pos_dat_begin Downto pos_dat_begin - 7) := data;
        End Loop;
        Return result;
    End Function;

    -------------------------------------------
    -- Set same the specified row of all digits
    -------------------------------------------
    Function clr_row(row_selector : RowSelectorType) Return DataStreamType Is
    Begin
        Return set_row(row_selector, "00000000");
    End Function;

    Constant REG_BCD_ENCODE      : RegType  := "1001";
    Constant D_BCD_ENCODE_NONE : DataType := "00000000";

    Constant REG_INTENSITY : RegType := "1010";
    Type IntensityType Is Array (0 To 15) Of DataType;
    Constant D_INTENSITY : IntensityType := (
        "00000000", "00000001", "00000010", "00000011", "00000100", "00000101", "00000110", "00000111",
        "00001000", "00001001", "00001010", "00001011", "00001100", "00001101", "00001110", "00001111"
    );

    ------------------------------------
    -- Intensity generator for digits --
    ------------------------------------

    Subtype DigitSelectorType Is std_logic_vector(19 Downto 0);
    Subtype IntensitySelectorType Is natural Range 0 To 15;
    Function set_intensity(digit_selectors    : DigitSelectorType;
                           intensity_selector : IntensitySelectorType) Return DataStreamType Is
        Variable result : DataStreamType;
        Variable pos_hdr_begin : integer;
        Variable pos_reg_begin : integer;
        Variable pos_dat_begin : integer;
    Begin
        For digit In DigitSelectorType'Range Loop
            pos_hdr_begin := (digit + 1) * 16 - 1;
            pos_reg_begin := pos_hdr_begin - 4;
            pos_dat_begin := pos_reg_begin - 4;
            result(pos_hdr_begin Downto pos_hdr_begin - 3) := HDR;
            If digit_selectors(digit) = '1' Then
                result(pos_reg_begin Downto pos_reg_begin - 3) := REG_INTENSITY;
                result(pos_dat_begin Downto pos_dat_begin - 7) := D_INTENSITY(intensity_selector);
            Else
                result(pos_reg_begin Downto pos_reg_begin - 3) := REG_NOP;
                result(pos_dat_begin Downto pos_dat_begin - 7) := D_NOP;
        End If;
        End Loop;
        Return result;
    End Function;


    Constant REG_SCAN          : RegType  := "1011";
    Constant D_SCAN_0xxxxxxx : DataType := "00000000";
    Constant D_SCAN_01xxxxxx : DataType := "00000001";
    Constant D_SCAN_012xxxxx : DataType := "00000010";
    Constant D_SCAN_0123xxxx : DataType := "00000011";
    Constant D_SCAN_01234xxx : DataType := "00000100";
    Constant D_SCAN_012345xx : DataType := "00000101";
    Constant D_SCAN_0123456x : DataType := "00000110";
    Constant D_SCAN_01234567 : DataType := "00000111";

    -- Make sure all digits are scanned (displayed)
    Constant SCAN_01234567 : DataStreamType :=
        HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 &
        HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 &
        HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 &
        HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 &
        HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567 & HDR & REG_SCAN & D_SCAN_01234567;

    -- Disable BCD encoding
    Constant BCD_ENCODE_NONE : DataStreamType :=
        HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE &
        HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE &
        HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE &
        HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE &
        HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE & HDR & REG_BCD_ENCODE & D_BCD_ENCODE_NONE;

    Constant REG_SHUT        : RegType  := "1100";
    Constant D_SHUT_DOWN   : DataType := "00000000";
    Constant D_SHUT_NORMAL : DataType := "00000001";

    -- Switch to the normal regime from possible shutdown mode
    Constant SHUT_NORMAL : DataStreamType :=
        HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL &
        HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL &
        HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL &
        HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL &
        HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL & HDR & REG_SHUT & D_SHUT_NORMAL;

    Constant REG_TEST   : RegType  := "1111";
    Constant D_TEST_0 : DataType := "00000000";
    Constant D_TEST_1 : DataType := "00000001";

    --------------------------
    -- Digit test generator --
    --------------------------
    Function test_digit(digit_selectors : DigitSelectorType) Return DataStreamType Is
        Variable result : DataStreamType;
        Variable pos_hdr_begin : integer;
        Variable pos_reg_begin : integer;
        Variable pos_dat_begin : integer;
    Begin
        For digit In DigitSelectorType'Range Loop
            pos_hdr_begin := (digit + 1) * 16 - 1;
            pos_reg_begin := pos_hdr_begin - 4;
            pos_dat_begin := pos_reg_begin - 4;
            result(pos_hdr_begin Downto pos_hdr_begin - 3) := HDR;
            result(pos_reg_begin Downto pos_reg_begin - 3) := REG_TEST;
            If digit_selectors(digit) = '1' Then
                result(pos_dat_begin Downto pos_dat_begin - 7) := D_TEST_1;
            Else
                result(pos_dat_begin Downto pos_dat_begin - 7) := D_TEST_0;
            End If;
        End Loop;
        Return result;
    End Function;

    Type TestsType Is Array (natural range <>) Of DataStreamType;
    Constant TESTS_1 : TestsType := (

        SHUT_NORMAL,
        SCAN_01234567,
        BCD_ENCODE_NONE,

        test_digit(B"0000_0000_0000_0000_0000"),
        test_digit(B"1111_1111_1111_1111_1111"),
        test_digit(B"0000_0000_0000_0000_0000"),
        test_digit(B"0000_0000_0000_0000_0001"),
        test_digit(B"0000_0000_0000_0000_0010"),
        test_digit(B"0000_0000_0000_0000_0100"),
        test_digit(B"0000_0000_0000_0000_1000"),
        test_digit(B"0000_0000_0000_0001_0000"),
        test_digit(B"0000_0000_0000_0010_0000"),
        test_digit(B"0000_0000_0000_0100_0000"),
        test_digit(B"0000_0000_0000_1000_0000"),
        test_digit(B"0000_0000_0001_0000_0000"),
        test_digit(B"0000_0000_0010_0000_0000"),
        test_digit(B"0000_0000_0100_0000_0000"),
        test_digit(B"0000_0000_1000_0000_0000"),
        test_digit(B"0000_0001_0000_0000_0000"),
        test_digit(B"0000_0010_0000_0000_0000"),
        test_digit(B"0000_0100_0000_0000_0000"),
        test_digit(B"0000_1000_0000_0000_0000"),
        test_digit(B"0001_0000_0000_0000_0000"),
        test_digit(B"0010_0000_0000_0000_0000"),
        test_digit(B"0100_0000_0000_0000_0000"),
        test_digit(B"1000_0000_0000_0000_0000"),
        test_digit(B"0100_0000_0000_0000_0000"),
        test_digit(B"0010_0000_0000_0000_0000"),
        test_digit(B"0001_0000_0000_0000_0000"),
        test_digit(B"0000_1000_0000_0000_0000"),
        test_digit(B"0000_0100_0000_0000_0000"),
        test_digit(B"0000_0010_0000_0000_0000"),
        test_digit(B"0000_0001_0000_0000_0000"),
        test_digit(B"0000_0000_1000_0000_0000"),
        test_digit(B"0000_0000_0100_0000_0000"),
        test_digit(B"0000_0000_0010_0000_0000"),
        test_digit(B"0000_0000_0001_0000_0000"),
        test_digit(B"0000_0000_0000_1000_0000"),
        test_digit(B"0000_0000_0000_0100_0000"),
        test_digit(B"0000_0000_0000_0010_0000"),
        test_digit(B"0000_0000_0000_0001_0000"),
        test_digit(B"0000_0000_0000_0000_1000"),
        test_digit(B"0000_0000_0000_0000_0100"),
        test_digit(B"0000_0000_0000_0000_0010"),
        test_digit(B"0000_0000_0000_0000_0001"),
        test_digit(B"0000_0000_0000_0000_0000"),

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, "01010101"),
        set_row(1, "10101010"),
        set_row(2, "01010101"),
        set_row(3, "10101010"),
        set_row(4, "01010101"),
        set_row(5, "10101010"),
        set_row(6, "01010101"),
        set_row(7, "10101010"),

        set_intensity(B"1111_1111_1111_1111_1111", 0),
        set_intensity(B"1111_1111_1111_1111_1111", 1),
        set_intensity(B"1111_1111_1111_1111_1111", 2),
        set_intensity(B"1111_1111_1111_1111_1111", 3),
        set_intensity(B"1111_1111_1111_1111_1111", 4),
        set_intensity(B"1111_1111_1111_1111_1111", 5),
        set_intensity(B"1111_1111_1111_1111_1111", 6),
        set_intensity(B"1111_1111_1111_1111_1111", 7),
        set_intensity(B"1111_1111_1111_1111_1111", 8),
        set_intensity(B"1111_1111_1111_1111_1111", 9),
        set_intensity(B"1111_1111_1111_1111_1111", 10),
        set_intensity(B"1111_1111_1111_1111_1111", 11),
        set_intensity(B"1111_1111_1111_1111_1111", 12),
        set_intensity(B"1111_1111_1111_1111_1111", 13),
        set_intensity(B"1111_1111_1111_1111_1111", 14),
        set_intensity(B"1111_1111_1111_1111_1111", 15),
        set_intensity(B"1111_1111_1111_1111_1111", 14),
        set_intensity(B"1111_1111_1111_1111_1111", 13),
        set_intensity(B"1111_1111_1111_1111_1111", 12),
        set_intensity(B"1111_1111_1111_1111_1111", 11),
        set_intensity(B"1111_1111_1111_1111_1111", 10),
        set_intensity(B"1111_1111_1111_1111_1111", 9),
        set_intensity(B"1111_1111_1111_1111_1111", 8),
        set_intensity(B"1111_1111_1111_1111_1111", 7),
        set_intensity(B"1111_1111_1111_1111_1111", 6),
        set_intensity(B"1111_1111_1111_1111_1111", 5),
        set_intensity(B"1111_1111_1111_1111_1111", 4),
        set_intensity(B"1111_1111_1111_1111_1111", 3),
        set_intensity(B"1111_1111_1111_1111_1111", 2),
        set_intensity(B"1111_1111_1111_1111_1111", 1),
        set_intensity(B"1111_1111_1111_1111_1111", 0),

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(0), 0)),
        set_row(1, symbol_row(DECIMAL(0), 1)),
        set_row(2, symbol_row(DECIMAL(0), 2)),
        set_row(3, symbol_row(DECIMAL(0), 3)),
        set_row(4, symbol_row(DECIMAL(0), 4)),
        set_row(5, symbol_row(DECIMAL(0), 5)),
        set_row(6, symbol_row(DECIMAL(0), 6)),
        set_row(7, symbol_row(DECIMAL(0), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(1), 0)),
        set_row(1, symbol_row(DECIMAL(1), 1)),
        set_row(2, symbol_row(DECIMAL(1), 2)),
        set_row(3, symbol_row(DECIMAL(1), 3)),
        set_row(4, symbol_row(DECIMAL(1), 4)),
        set_row(5, symbol_row(DECIMAL(1), 5)),
        set_row(6, symbol_row(DECIMAL(1), 6)),
        set_row(7, symbol_row(DECIMAL(1), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(2), 0)),
        set_row(1, symbol_row(DECIMAL(2), 1)),
        set_row(2, symbol_row(DECIMAL(2), 2)),
        set_row(3, symbol_row(DECIMAL(2), 3)),
        set_row(4, symbol_row(DECIMAL(2), 4)),
        set_row(5, symbol_row(DECIMAL(2), 5)),
        set_row(6, symbol_row(DECIMAL(2), 6)),
        set_row(7, symbol_row(DECIMAL(2), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(3), 0)),
        set_row(1, symbol_row(DECIMAL(3), 1)),
        set_row(2, symbol_row(DECIMAL(3), 2)),
        set_row(3, symbol_row(DECIMAL(3), 3)),
        set_row(4, symbol_row(DECIMAL(3), 4)),
        set_row(5, symbol_row(DECIMAL(3), 5)),
        set_row(6, symbol_row(DECIMAL(3), 6)),
        set_row(7, symbol_row(DECIMAL(3), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(4), 0)),
        set_row(1, symbol_row(DECIMAL(4), 1)),
        set_row(2, symbol_row(DECIMAL(4), 2)),
        set_row(3, symbol_row(DECIMAL(4), 3)),
        set_row(4, symbol_row(DECIMAL(4), 4)),
        set_row(5, symbol_row(DECIMAL(4), 5)),
        set_row(6, symbol_row(DECIMAL(4), 6)),
        set_row(7, symbol_row(DECIMAL(4), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(5), 0)),
        set_row(1, symbol_row(DECIMAL(5), 1)),
        set_row(2, symbol_row(DECIMAL(5), 2)),
        set_row(3, symbol_row(DECIMAL(5), 3)),
        set_row(4, symbol_row(DECIMAL(5), 4)),
        set_row(5, symbol_row(DECIMAL(5), 5)),
        set_row(6, symbol_row(DECIMAL(5), 6)),
        set_row(7, symbol_row(DECIMAL(5), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(6), 0)),
        set_row(1, symbol_row(DECIMAL(6), 1)),
        set_row(2, symbol_row(DECIMAL(6), 2)),
        set_row(3, symbol_row(DECIMAL(6), 3)),
        set_row(4, symbol_row(DECIMAL(6), 4)),
        set_row(5, symbol_row(DECIMAL(6), 5)),
        set_row(6, symbol_row(DECIMAL(6), 6)),
        set_row(7, symbol_row(DECIMAL(6), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(7), 0)),
        set_row(1, symbol_row(DECIMAL(7), 1)),
        set_row(2, symbol_row(DECIMAL(7), 2)),
        set_row(3, symbol_row(DECIMAL(7), 3)),
        set_row(4, symbol_row(DECIMAL(7), 4)),
        set_row(5, symbol_row(DECIMAL(7), 5)),
        set_row(6, symbol_row(DECIMAL(7), 6)),
        set_row(7, symbol_row(DECIMAL(7), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(8), 0)),
        set_row(1, symbol_row(DECIMAL(8), 1)),
        set_row(2, symbol_row(DECIMAL(8), 2)),
        set_row(3, symbol_row(DECIMAL(8), 3)),
        set_row(4, symbol_row(DECIMAL(8), 4)),
        set_row(5, symbol_row(DECIMAL(8), 5)),
        set_row(6, symbol_row(DECIMAL(8), 6)),
        set_row(7, symbol_row(DECIMAL(8), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP,

        clr_row(7), clr_row(6), clr_row(5), clr_row(4), clr_row(3), clr_row(2), clr_row(1), clr_row(0),

        set_row(0, symbol_row(DECIMAL(9), 0)),
        set_row(1, symbol_row(DECIMAL(9), 1)),
        set_row(2, symbol_row(DECIMAL(9), 2)),
        set_row(3, symbol_row(DECIMAL(9), 3)),
        set_row(4, symbol_row(DECIMAL(9), 4)),
        set_row(5, symbol_row(DECIMAL(9), 5)),
        set_row(6, symbol_row(DECIMAL(9), 6)),
        set_row(7, symbol_row(DECIMAL(9), 7)),

        NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP, NOP
    );
    Signal data : DataStreamType;

    -- Rotary encoder driving the level meter

    Constant METER_WIDTH : positive := positive(ceil(log2(real(10**DIGITS))));

    Constant METERED_VAL_0 : unsigned(METER_WIDTH - 1 Downto 0) := to_unsigned(10,   METER_WIDTH);
    Constant METERED_VAL_1 : unsigned(METER_WIDTH - 1 Downto 0) := to_unsigned(100,  METER_WIDTH);
    Constant METERED_VAL_2 : unsigned(METER_WIDTH - 1 Downto 0) := to_unsigned(1000, METER_WIDTH);
    Constant METERED_VAL_3 : unsigned(METER_WIDTH - 1 Downto 0) := to_unsigned(2000, METER_WIDTH);

    Signal metered_value     : std_logic_vector(METER_WIDTH - 1 Downto 0) := (Others => '0');
    Signal metered_bcd_value : std_logic_vector(DIGITS * 4 - 1 Downto 0) := (Others => '0');
    Signal counter_clk       : std_logic;

    Signal metered_value_0 : unsigned(METER_WIDTH - 1 Downto 0) := (Others => '0');
    Signal metered_value_1 : unsigned(METER_WIDTH - 1 Downto 0) := (Others => '0');
    Signal metered_value_2 : unsigned(METER_WIDTH - 1 Downto 0) := (Others => '0');
    Signal metered_value_3 : unsigned(METER_WIDTH - 1 Downto 0) := (Others => '0');

    Signal TESTS_2 : TestsType := (
        SHUT_NORMAL,
        SHUT_NORMAL,
        SCAN_01234567,
        SCAN_01234567,
        BCD_ENCODE_NONE,
        BCD_ENCODE_NONE,
        set_intensity(B"1111_1111_1111_1111_1111", 15),
        set_intensity(B"1111_1111_1111_1111_1111", 15),
        set_row(0, symbol_row(DECIMAL(0), 0)),
        set_row(1, symbol_row(DECIMAL(0), 1)),
        set_row(2, symbol_row(DECIMAL(0), 2)),
        set_row(3, symbol_row(DECIMAL(0), 3)),
        set_row(4, symbol_row(DECIMAL(0), 4)),
        set_row(5, symbol_row(DECIMAL(0), 5)),
        set_row(6, symbol_row(DECIMAL(0), 6)),
        set_row(7, symbol_row(DECIMAL(0), 7))
    );

    -- Debounced push buttons on the rotary encoder driving the level meter.
    Signal rencoder_btn : std_logic_vector(0 To DIGITS - 1);

    Component c_addsub_0
        Port(A   : In unsigned(METER_WIDTH - 1 Downto 0);
             B   : In unsigned(METER_WIDTH - 1 Downto 0);
             CLK : In std_logic;
             S   : Out unsigned(METER_WIDTH - 1 Downto 0)
        );
    End Component;

Begin

    -- Running sums
    adder_0 : c_addsub_0
        Port Map(A   => unsigned(metered_value),
                 B   => METERED_VAL_0,
                 CLK => clk,
                 S   => metered_value_0);

    adder_1 : c_addsub_0
        Port Map(A   => unsigned(metered_value),
                 B   => METERED_VAL_1,
                 CLK => clk,
                 S   => metered_value_1);

    adder_2 : c_addsub_0
        Port Map(A   => unsigned(metered_value),
                 B   => METERED_VAL_2,
                 CLK => clk,
                 S   => metered_value_2);

    adder_3 : c_addsub_0
        Port Map(A   => unsigned(metered_value),
                 B   => METERED_VAL_3,
                 CLK => clk,
                 S   => metered_value_3);
        
    -- Debouncers for the eeset button and the rotary encoder buttons.
    rst_button_debouncer : Entity work.debouncer
        Generic Map(CLK_PERIODS => FREQ_RENCODER_CLK_PERIODS)
        Port    Map(i_clk => clk,
                    i_btn => rst_btn,
                    o_btn => rst);

    generate_rencoder_buttons : For idx In 0 To DIGITS - 1 Generate
        button_debouncer : Entity work.debouncer
            Generic Map(CLK_PERIODS => FREQ_RENCODER_CLK_PERIODS)
            Port    Map(i_clk => clk,
                        i_btn => Not g_rencoder_p(idx),
                        o_btn => rencoder_btn(idx));
    End Generate generate_rencoder_buttons;

    g_rencoder_left  <= rencoder_btn(0);
    g_rencoder_right <= rencoder_btn(1);

    -- LED display update process keeps selecting the content of the framebuffer
    -- stream by stream and updating the data register. The register is pushed
    -- next to the LED matrix via SPI.
    display_update_process : Process (spi_drive_clk, rst) Is
        Alias TESTS : TestsType Is TESTS_2;
        Constant MAX_CYCLES : natural := FREQ_SPI_DRIVE_CLK / FREQ_DISPLEY_UPDATE;
        Variable num_cycles : natural := 0;
        Variable test_idx   : natural := TESTS'Left;
    Begin
        If rst Then
            num_cycles := 0;
            test_idx := TESTS'Left;
            start <= '0';
        Else
            If rising_edge(spi_drive_clk) Then
                If Not busy Then
                    num_cycles := num_cycles + 1;
                    If num_cycles = MAX_CYCLES Then
                        num_cycles := 0;
                        data <= TESTS(test_idx);
                        If test_idx = TESTS'Right Then
                            test_idx := TESTS'Left;
                        Else
                            test_idx := test_idx + 1;
                        End If;
                        start <= '1';
                    Else
                        start <= '0';
                    End If;
                End If;
            End If;    
        End If;
    End Process display_update_process;

    -- Clock divider to make the desired clock driving the module
    clock_driver :
        Entity work.clock_div
            Generic Map(N => FREQ_CLK / FREQ_SPI_DRIVE_CLK)
            Port    Map(i_rst => rst,
                        i_clk => clk,
                        o_clk => spi_drive_clk);

    -- A driver for the SPI signals generator
    max7219_driver :
        Entity work.spi_max7219_synt
            Generic Map(WIDTH => DataStreamType'Length)
            Port Map(i_rst        => rst,
                     i_clk        => spi_drive_clk,
                     i_start      => start,
                     i_data       => data,
                     o_busy       => busy,
                     o_spi_clk    => g_spi_clk,
                     o_spi_load   => spi_load,
                     o_spi_din    => g_spi_din,
                     o_diag_state => diag_state);

    g_spi_load <= spi_load;
    g_div_clk  <= spi_drive_clk;

    ---------------------------------------------------------------------------------
    -- Temporarily disabled to allow runing the clock-driven increment of the metered
    -- value instead of using knobs.
    --
    -- rencoder_driver :
    --     Entity work.meter_n
    --         Generic Map(CLK_PERIODS => FREQ_RENCODER_CLK_PERIODS,
    --                     DIGITS => DIGITS,
    --                     METER_WIDTH => METER_WIDTH)
    --         Port    Map(i_clk   => clk,
    --                     i_a     => g_rencoder_a(0 To DIGITS-1),
    --                     i_b     => g_rencoder_b(0 To DIGITS-1),
    --                     o_value => metered_value);

    ----------------------------------------------------------------------------------
    -- This is just a test for how the encoder works. The output is sent to the output
    -- ports of the FPGA.
    -- rencoder_driver_4 :
    --     Entity work.encoder
    --         Generic Map(CLK_PERIODS => FREQ_RENCODER_CLK_PERIODS)
    --         Port    Map(i_clk   => clk,
    --                     i_a     => g_rencoder_a(4),
    --                     i_b     => g_rencoder_b(4),
    --                     o_left  => g_rencoder_left,
    --                     o_right => g_rencoder_right);

    ------------------------------------------------------------------------------------
    -- Clock divider to make the clock driving a process incrementing the metered value.
    -- This is just a test for the display.

    counter_clock_driver :
        Entity work.clock_div
            Generic Map(N => FREQ_CLK / FREQ_COUNTER_CLK)
            Port    Map(i_rst => rst,
                        i_clk => clk,
                        o_clk => counter_clk);

    counter_increment_process : Process (counter_clk, rst, rencoder_btn) Is
    Begin
        If rst Then
            metered_value <= (Others => '0');
        ElsIf rencoder_btn(0) Then
            metered_value <= std_logic_vector(metered_value_0);
        ElsIf rencoder_btn(1) Then
            metered_value <= std_logic_vector(metered_value_1);
        ElsIf rencoder_btn(2) Then
            metered_value <= std_logic_vector(metered_value_2);
        ElsIf rencoder_btn(3) Then
            metered_value <= std_logic_vector(metered_value_3);
        ElsIf rising_edge(counter_clk) Then
            metered_value <= metered_value + '1';
        End If;
    End Process counter_increment_process;

    decoder_bin2bcd : Entity work.decod_bin2bcd_para
    Generic Map(INPUT_WIDTH    => METER_WIDTH,
                DECIMAL_DIGITS => DIGITS)
    Port    Map(bin => metered_value,
                bcd => metered_bcd_value);

    ----------------------------------------------------------------------------------
    -- This process updates the BCD number on the display each time the value changes.
    --
    -- COMMENTS/QUESTIONS:
    -- a) The process is triggered by changes in the BCD value, which seems to work fine
    -- b) However the processs updates the framebuffer of the display using operator <=
    -- c) Does this mean that the framebuffer is allocated in the block memory rather than
    --    using triiggers? 

    test_update: For row In 0 To 7 Generate
        test_update_process : Process (metered_bcd_value) Is
            Variable idx0 : integer;
            Variable idx1 : integer;
            Variable idx2 : integer;
            Variable idx3 : integer;
        Begin
            idx0 := to_integer(unsigned(metered_bcd_value( 3 Downto  0)));
            idx1 := to_integer(unsigned(metered_bcd_value( 7 Downto  4)));
            idx2 := to_integer(unsigned(metered_bcd_value(11 Downto  8)));
            idx3 := to_integer(unsigned(metered_bcd_value(15 Downto 12)));
            TESTS_2(8 + row) <=
                HDR & REG_ROW(row) & symbol_row(DECIMAL(idx0), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx1), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx2), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx3), row) &
                HDR & REG_ROW(row) & symbol_row(DECIMAL(idx0), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx1), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx2), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx3), row) &
                HDR & REG_ROW(row) & symbol_row(DECIMAL(idx0), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx1), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx2), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx3), row) &
                HDR & REG_ROW(row) & symbol_row(DECIMAL(idx0), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx1), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx2), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx3), row) &
                HDR & REG_ROW(row) & symbol_row(DECIMAL(idx0), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx1), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx2), row) & HDR & REG_ROW(row) & symbol_row(DECIMAL(idx3), row);
        End Process test_update_process;
    End Generate test_update;

End Architecture Rtl;
