fb[36][13] <= 1'b1;
fb[36][15] <= 1'b1;
fb[36][17] <= 1'b1;
fb[35][9] <= 1'b1;
fb[35][21] <= 1'b1;
fb[34][7] <= 1'b1;
fb[34][23] <= 1'b1;
fb[32][5] <= 1'b1;
fb[32][25] <= 1'b1;
fb[31][4] <= 1'b1;
fb[31][26] <= 1'b1;
fb[29][3] <= 1'b1;
fb[29][27] <= 1'b1;
fb[25][2] <= 1'b1;
fb[25][28] <= 1'b1;
fb[23][2] <= 1'b1;
fb[23][28] <= 1'b1;
fb[21][2] <= 1'b1;
fb[21][28] <= 1'b1;
fb[17][3] <= 1'b1;
fb[17][27] <= 1'b1;
fb[15][4] <= 1'b1;
fb[15][26] <= 1'b1;
fb[14][5] <= 1'b1;
fb[14][25] <= 1'b1;
fb[12][7] <= 1'b1;
fb[12][23] <= 1'b1;
fb[11][9] <= 1'b1;
fb[11][21] <= 1'b1;
fb[10][13] <= 1'b1;
fb[10][15] <= 1'b1;
fb[10][17] <= 1'b1;
fb[6][14] <= 1'b1;
fb[6][16] <= 1'b1;
fb[6][17] <= 1'b1;
fb[6][18] <= 1'b1;
fb[6][19] <= 1'b1;
fb[6][20] <= 1'b1;
fb[5][14] <= 1'b1;
fb[5][20] <= 1'b1;
fb[4][14] <= 1'b1;
fb[4][20] <= 1'b1;
fb[3][14] <= 1'b1;
fb[3][16] <= 1'b1;
fb[3][17] <= 1'b1;
fb[3][18] <= 1'b1;
fb[3][19] <= 1'b1;
fb[3][20] <= 1'b1;
fb[2][14] <= 1'b1;
fb[2][20] <= 1'b1;
fb[1][14] <= 1'b1;
fb[1][20] <= 1'b1;
fb[0][14] <= 1'b1;
fb[0][16] <= 1'b1;
fb[0][17] <= 1'b1;
fb[0][18] <= 1'b1;
fb[0][19] <= 1'b1;
fb[0][20] <= 1'b1;
