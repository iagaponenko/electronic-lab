fb[34][13] <= 1'b1;
fb[34][15] <= 1'b1;
fb[34][17] <= 1'b1;
fb[33][10] <= 1'b1;
fb[33][20] <= 1'b1;
fb[32][8] <= 1'b1;
fb[32][22] <= 1'b1;
fb[31][7] <= 1'b1;
fb[31][23] <= 1'b1;
fb[30][6] <= 1'b1;
fb[30][24] <= 1'b1;
fb[28][5] <= 1'b1;
fb[28][25] <= 1'b1;
fb[25][4] <= 1'b1;
fb[25][26] <= 1'b1;
fb[23][4] <= 1'b1;
fb[23][26] <= 1'b1;
fb[21][4] <= 1'b1;
fb[21][26] <= 1'b1;
fb[18][5] <= 1'b1;
fb[18][25] <= 1'b1;
fb[16][6] <= 1'b1;
fb[16][24] <= 1'b1;
fb[15][7] <= 1'b1;
fb[15][23] <= 1'b1;
fb[14][8] <= 1'b1;
fb[14][22] <= 1'b1;
fb[13][10] <= 1'b1;
fb[13][20] <= 1'b1;
fb[12][13] <= 1'b1;
fb[12][15] <= 1'b1;
fb[12][17] <= 1'b1;
fb[6][14] <= 1'b1;
fb[6][20] <= 1'b1;
fb[5][14] <= 1'b1;
fb[5][20] <= 1'b1;
fb[4][14] <= 1'b1;
fb[4][20] <= 1'b1;
fb[3][14] <= 1'b1;
fb[3][20] <= 1'b1;
fb[2][14] <= 1'b1;
fb[2][20] <= 1'b1;
fb[1][14] <= 1'b1;
fb[1][20] <= 1'b1;
fb[0][14] <= 1'b1;
fb[0][20] <= 1'b1;
