-- Implement an SPI-like serializer for MAX7219.
-- The syntesizable version in which each SPI clock period is 3 times
-- longer than the input clock.
--
-- https://www.sparkfun.com/datasheets/Components/General/COM-09622-MAX7219-MAX7221.pdf

Library ieee;
Use ieee.std_logic_1164.All;
Use ieee.numeric_std.All;
Use ieee.math_real.All;

Entity spi_max7219_synt Is
    Port (
        -- Management interface
        i_rst        : In  std_logic;
        i_clk        : In  std_logic;
        i_start      : In  std_logic;
        i_data       : In  std_logic_vector(15 Downto 0);
        o_busy       : Out std_logic;
        -- SPI signals generated by the entity
        o_spi_clk    : Out std_logic;
        o_spi_load   : Out std_logic;
        o_spi_din    : Out std_logic;
        -- Diagnostics
        o_diag_state : Out std_logic_vector(1 Downto 0)
    );
End Entity spi_max7219_synt;

Architecture Rtl Of spi_max7219_synt Is
    Type ProcessingState Is (IDLE, DATA_IN, CLOCK_RISE, CLOCK_FALL);
    Signal state : ProcessingState;
Begin
    bcd_compute_process : Process (i_clk, i_rst) Is
        Variable index : integer Range 0 To 15;
    Begin
        If i_rst Then
            state <= IDLE;
        ElsIf rising_edge(i_clk) Then
            Case state Is
                When IDLE =>
                    o_spi_clk  <= '0';
                    o_spi_load <= '0';
                    o_spi_din  <= 'X';
                    If i_start Then
                        index := 15;
                        state <= DATA_IN;
                    End If;
                When DATA_IN =>
                    o_spi_din <= i_data(index);
                    state <= CLOCK_RISE;
                When CLOCK_RISE =>
                    o_spi_clk <= '1';
--                     If index = 0 Then
--                         o_spi_load <= '1';
--                     End If;
                    state <= CLOCK_FALL;
                When CLOCK_FALL =>
                    o_spi_clk <= '0';
                    If index = 0 Then
                        o_spi_load <= '1';
                        state <= IDLE;
                    Else
                        index := index - 1;
                        state <= DATA_IN;
                    End If;
                When Others =>
                    state <= IDLE;
            End Case;
        End If;
    End Process bcd_compute_process;

    -- Device "o_busy" is set during when the last request is still being processed.
    -- The "i_start" command will be ignored in this state.
    o_busy <= '0' When state = IDLE       Else
              '1' When state = DATA_IN    Else
              '1' When state = CLOCK_RISE Else
              '1' When state = CLOCK_FALL Else
              'X';

    -- Diagnostic signals
    o_diag_state <= "00" When state = IDLE       Else
                    "01" When state = DATA_IN    Else
                    "10" When state = CLOCK_RISE Else
                    "11" When state = CLOCK_FALL Else
                    "XX";

End Architecture Rtl;

