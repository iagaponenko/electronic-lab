fb[25][14] <= 1'b0;
fb[25][15] <= 1'b0;
fb[25][16] <= 1'b0;
fb[24][13] <= 1'b0;
fb[24][17] <= 1'b0;
fb[23][13] <= 1'b0;
fb[23][17] <= 1'b0;
fb[22][13] <= 1'b0;
fb[22][17] <= 1'b0;
fb[21][14] <= 1'b0;
fb[21][15] <= 1'b0;
fb[21][16] <= 1'b0;
fb[6][10] <= 1'b0;
fb[6][11] <= 1'b0;
fb[6][12] <= 1'b0;
fb[6][13] <= 1'b0;
fb[6][14] <= 1'b0;
fb[6][16] <= 1'b0;
fb[6][17] <= 1'b0;
fb[6][18] <= 1'b0;
fb[6][19] <= 1'b0;
fb[6][20] <= 1'b0;
fb[5][10] <= 1'b0;
fb[5][14] <= 1'b0;
fb[5][20] <= 1'b0;
fb[4][10] <= 1'b0;
fb[4][14] <= 1'b0;
fb[4][20] <= 1'b0;
fb[3][10] <= 1'b0;
fb[3][14] <= 1'b0;
fb[3][16] <= 1'b0;
fb[3][17] <= 1'b0;
fb[3][18] <= 1'b0;
fb[3][19] <= 1'b0;
fb[3][20] <= 1'b0;
fb[2][10] <= 1'b0;
fb[2][14] <= 1'b0;
fb[2][16] <= 1'b0;
fb[1][10] <= 1'b0;
fb[1][14] <= 1'b0;
fb[1][16] <= 1'b0;
fb[0][10] <= 1'b0;
fb[0][11] <= 1'b0;
fb[0][12] <= 1'b0;
fb[0][13] <= 1'b0;
fb[0][14] <= 1'b0;
fb[0][16] <= 1'b0;
fb[0][17] <= 1'b0;
fb[0][18] <= 1'b0;
fb[0][19] <= 1'b0;
fb[0][20] <= 1'b0;
