fb[39][12] <= 1'b1;
fb[39][15] <= 1'b1;
fb[39][18] <= 1'b1;
fb[38][9] <= 1'b1;
fb[38][21] <= 1'b1;
fb[37][7] <= 1'b1;
fb[37][23] <= 1'b1;
fb[35][4] <= 1'b1;
fb[35][26] <= 1'b1;
fb[33][2] <= 1'b1;
fb[33][28] <= 1'b1;
fb[31][1] <= 1'b1;
fb[31][29] <= 1'b1;
fb[29][0] <= 1'b1;
fb[29][30] <= 1'b1;
fb[26][31] <= 1'b1;
fb[23][31] <= 1'b1;
fb[20][31] <= 1'b1;
fb[17][0] <= 1'b1;
fb[17][30] <= 1'b1;
fb[15][1] <= 1'b1;
fb[15][29] <= 1'b1;
fb[13][2] <= 1'b1;
fb[13][28] <= 1'b1;
fb[11][4] <= 1'b1;
fb[11][26] <= 1'b1;
fb[9][7] <= 1'b1;
fb[9][23] <= 1'b1;
fb[8][9] <= 1'b1;
fb[8][21] <= 1'b1;
fb[6][14] <= 1'b1;
fb[6][16] <= 1'b1;
fb[6][17] <= 1'b1;
fb[6][18] <= 1'b1;
fb[6][19] <= 1'b1;
fb[6][20] <= 1'b1;
fb[5][14] <= 1'b1;
fb[5][16] <= 1'b1;
fb[4][14] <= 1'b1;
fb[4][16] <= 1'b1;
fb[3][14] <= 1'b1;
fb[3][16] <= 1'b1;
fb[3][17] <= 1'b1;
fb[3][18] <= 1'b1;
fb[3][19] <= 1'b1;
fb[3][20] <= 1'b1;
fb[2][14] <= 1'b1;
fb[2][16] <= 1'b1;
fb[2][20] <= 1'b1;
fb[1][14] <= 1'b1;
fb[1][16] <= 1'b1;
fb[1][20] <= 1'b1;
fb[0][14] <= 1'b1;
fb[0][16] <= 1'b1;
fb[0][17] <= 1'b1;
fb[0][18] <= 1'b1;
fb[0][19] <= 1'b1;
fb[0][20] <= 1'b1;
