fb[31][14] <= 1'b0;
fb[31][16] <= 1'b0;
fb[30][12] <= 1'b0;
fb[30][18] <= 1'b0;
fb[29][10] <= 1'b0;
fb[29][20] <= 1'b0;
fb[28][9] <= 1'b0;
fb[28][21] <= 1'b0;
fb[26][8] <= 1'b0;
fb[26][22] <= 1'b0;
fb[24][7] <= 1'b0;
fb[24][23] <= 1'b0;
fb[22][7] <= 1'b0;
fb[22][23] <= 1'b0;
fb[20][8] <= 1'b0;
fb[20][22] <= 1'b0;
fb[18][9] <= 1'b0;
fb[18][21] <= 1'b0;
fb[17][10] <= 1'b0;
fb[17][20] <= 1'b0;
fb[16][12] <= 1'b0;
fb[16][18] <= 1'b0;
fb[15][14] <= 1'b0;
fb[15][16] <= 1'b0;
fb[6][10] <= 1'b0;
fb[6][11] <= 1'b0;
fb[6][12] <= 1'b0;
fb[6][13] <= 1'b0;
fb[6][14] <= 1'b0;
fb[6][16] <= 1'b0;
fb[6][17] <= 1'b0;
fb[6][18] <= 1'b0;
fb[6][19] <= 1'b0;
fb[6][20] <= 1'b0;
fb[5][10] <= 1'b0;
fb[5][14] <= 1'b0;
fb[5][16] <= 1'b0;
fb[5][20] <= 1'b0;
fb[4][10] <= 1'b0;
fb[4][14] <= 1'b0;
fb[4][16] <= 1'b0;
fb[4][20] <= 1'b0;
fb[3][10] <= 1'b0;
fb[3][14] <= 1'b0;
fb[3][16] <= 1'b0;
fb[3][17] <= 1'b0;
fb[3][18] <= 1'b0;
fb[3][19] <= 1'b0;
fb[3][20] <= 1'b0;
fb[2][10] <= 1'b0;
fb[2][14] <= 1'b0;
fb[2][16] <= 1'b0;
fb[2][20] <= 1'b0;
fb[1][10] <= 1'b0;
fb[1][14] <= 1'b0;
fb[1][16] <= 1'b0;
fb[1][20] <= 1'b0;
fb[0][10] <= 1'b0;
fb[0][11] <= 1'b0;
fb[0][12] <= 1'b0;
fb[0][13] <= 1'b0;
fb[0][14] <= 1'b0;
fb[0][16] <= 1'b0;
fb[0][17] <= 1'b0;
fb[0][18] <= 1'b0;
fb[0][19] <= 1'b0;
fb[0][20] <= 1'b0;
