fb[35][13] <= 1'b0;
fb[35][15] <= 1'b0;
fb[35][17] <= 1'b0;
fb[34][10] <= 1'b0;
fb[34][20] <= 1'b0;
fb[33][8] <= 1'b0;
fb[33][22] <= 1'b0;
fb[31][6] <= 1'b0;
fb[31][24] <= 1'b0;
fb[30][5] <= 1'b0;
fb[30][25] <= 1'b0;
fb[28][4] <= 1'b0;
fb[28][26] <= 1'b0;
fb[25][3] <= 1'b0;
fb[25][27] <= 1'b0;
fb[23][3] <= 1'b0;
fb[23][27] <= 1'b0;
fb[21][3] <= 1'b0;
fb[21][27] <= 1'b0;
fb[18][4] <= 1'b0;
fb[18][26] <= 1'b0;
fb[16][5] <= 1'b0;
fb[16][25] <= 1'b0;
fb[15][6] <= 1'b0;
fb[15][24] <= 1'b0;
fb[13][8] <= 1'b0;
fb[13][22] <= 1'b0;
fb[12][10] <= 1'b0;
fb[12][20] <= 1'b0;
fb[11][13] <= 1'b0;
fb[11][15] <= 1'b0;
fb[11][17] <= 1'b0;
fb[6][14] <= 1'b0;
fb[6][16] <= 1'b0;
fb[6][17] <= 1'b0;
fb[6][18] <= 1'b0;
fb[6][19] <= 1'b0;
fb[6][20] <= 1'b0;
fb[5][14] <= 1'b0;
fb[5][20] <= 1'b0;
fb[4][14] <= 1'b0;
fb[4][20] <= 1'b0;
fb[3][14] <= 1'b0;
fb[3][16] <= 1'b0;
fb[3][17] <= 1'b0;
fb[3][18] <= 1'b0;
fb[3][19] <= 1'b0;
fb[3][20] <= 1'b0;
fb[2][14] <= 1'b0;
fb[2][16] <= 1'b0;
fb[1][14] <= 1'b0;
fb[1][16] <= 1'b0;
fb[0][14] <= 1'b0;
fb[0][16] <= 1'b0;
fb[0][17] <= 1'b0;
fb[0][18] <= 1'b0;
fb[0][19] <= 1'b0;
fb[0][20] <= 1'b0;
