fb[32][14] <= 1'b0;
fb[32][16] <= 1'b0;
fb[31][11] <= 1'b0;
fb[31][19] <= 1'b0;
fb[30][9] <= 1'b0;
fb[30][21] <= 1'b0;
fb[29][8] <= 1'b0;
fb[29][22] <= 1'b0;
fb[27][7] <= 1'b0;
fb[27][23] <= 1'b0;
fb[24][6] <= 1'b0;
fb[24][24] <= 1'b0;
fb[22][6] <= 1'b0;
fb[22][24] <= 1'b0;
fb[19][7] <= 1'b0;
fb[19][23] <= 1'b0;
fb[17][8] <= 1'b0;
fb[17][22] <= 1'b0;
fb[16][9] <= 1'b0;
fb[16][21] <= 1'b0;
fb[15][11] <= 1'b0;
fb[15][19] <= 1'b0;
fb[14][14] <= 1'b0;
fb[14][16] <= 1'b0;
fb[6][10] <= 1'b0;
fb[6][11] <= 1'b0;
fb[6][12] <= 1'b0;
fb[6][13] <= 1'b0;
fb[6][14] <= 1'b0;
fb[6][16] <= 1'b0;
fb[6][17] <= 1'b0;
fb[6][18] <= 1'b0;
fb[6][19] <= 1'b0;
fb[6][20] <= 1'b0;
fb[5][10] <= 1'b0;
fb[5][14] <= 1'b0;
fb[5][16] <= 1'b0;
fb[5][20] <= 1'b0;
fb[4][10] <= 1'b0;
fb[4][14] <= 1'b0;
fb[4][16] <= 1'b0;
fb[4][20] <= 1'b0;
fb[3][10] <= 1'b0;
fb[3][14] <= 1'b0;
fb[3][16] <= 1'b0;
fb[3][17] <= 1'b0;
fb[3][18] <= 1'b0;
fb[3][19] <= 1'b0;
fb[3][20] <= 1'b0;
fb[2][10] <= 1'b0;
fb[2][14] <= 1'b0;
fb[2][20] <= 1'b0;
fb[1][10] <= 1'b0;
fb[1][14] <= 1'b0;
fb[1][20] <= 1'b0;
fb[0][10] <= 1'b0;
fb[0][11] <= 1'b0;
fb[0][12] <= 1'b0;
fb[0][13] <= 1'b0;
fb[0][14] <= 1'b0;
fb[0][20] <= 1'b0;
